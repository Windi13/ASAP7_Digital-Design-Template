module counter_board (clock_i,
    enable_i,
    reset_n_i,
    counter_value_o);
 input clock_i;
 input enable_i;
 input reset_n_i;
 output [3:0] counter_value_o;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire clknet_0_clock_i;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net1;
 wire net2;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_1_0__leaf_clock_i;
 wire clknet_1_1__leaf_clock_i;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;

 INVx1_ASAP7_75t_R _19_ (.A(_00_),
    .Y(net6));
 INVx2_ASAP7_75t_R _20_ (.A(_01_),
    .Y(net5));
 INVx2_ASAP7_75t_R _21_ (.A(_02_),
    .Y(net4));
 INVx2_ASAP7_75t_R _22_ (.A(_03_),
    .Y(net3));
 INVx2_ASAP7_75t_R _23_ (.A(net2),
    .Y(_10_));
 OR3x1_ASAP7_75t_R _24_ (.A(_04_),
    .B(_01_),
    .C(_00_),
    .Y(_11_));
 AND3x1_ASAP7_75t_R _25_ (.A(_11_),
    .B(net2),
    .C(net14),
    .Y(_12_));
 AO21x1_ASAP7_75t_R _26_ (.A1(net21),
    .A2(_10_),
    .B(_12_),
    .Y(_06_));
 NAND2x1_ASAP7_75t_R _27_ (.A(net2),
    .B(_05_),
    .Y(_13_));
 OA21x2_ASAP7_75t_R _28_ (.A1(net25),
    .A2(net2),
    .B(_13_),
    .Y(_07_));
 NOR2x2_ASAP7_75t_R _29_ (.A(net11),
    .B(_10_),
    .Y(_14_));
 XNOR2x1_ASAP7_75t_R _30_ (.B(_14_),
    .Y(_08_),
    .A(net22));
 OR4x1_ASAP7_75t_R _31_ (.A(net23),
    .B(net15),
    .C(net14),
    .D(_10_),
    .Y(_15_));
 OAI21x1_ASAP7_75t_R _32_ (.A1(net16),
    .A2(net13),
    .B(net12),
    .Y(_16_));
 AND4x1_ASAP7_75t_R _33_ (.A(_16_),
    .B(net5),
    .C(net2),
    .D(net6),
    .Y(_17_));
 AOI21x1_ASAP7_75t_R _34_ (.A1(_00_),
    .A2(_15_),
    .B(_17_),
    .Y(_09_));
 HAxp5_ASAP7_75t_R _35_ (.A(net4),
    .B(net3),
    .CON(_04_),
    .SN(_05_));
 BUFx2_ASAP7_75t_R clkbuf_0_clock_i (.A(clock_i),
    .Y(clknet_0_clock_i));
 DFFASRHQNx1_ASAP7_75t_R \counter_0.n20_q[0]$_DFFE_PN0P_  (.CLK(clknet_1_0__leaf_clock_i),
    .D(_06_),
    .QN(_03_),
    .RESETN(net7),
    .SETN(net1));
 DFFASRHQNx1_ASAP7_75t_R \counter_0.n20_q[1]$_DFFE_PN0P_  (.CLK(clknet_1_1__leaf_clock_i),
    .D(_07_),
    .QN(_02_),
    .RESETN(net8),
    .SETN(net1));
 DFFASRHQNx1_ASAP7_75t_R \counter_0.n20_q[2]$_DFFE_PN0P_  (.CLK(clknet_1_0__leaf_clock_i),
    .D(_08_),
    .QN(_01_),
    .RESETN(net9),
    .SETN(net1));
 DFFASRHQNx1_ASAP7_75t_R \counter_0.n20_q[3]$_DFFE_PN0P_  (.CLK(clknet_1_1__leaf_clock_i),
    .D(_09_),
    .QN(_00_),
    .RESETN(net10),
    .SETN(net1));
 BUFx2_ASAP7_75t_R hold1 (.A(net24),
    .Y(net1));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_57 ();
 BUFx2_ASAP7_75t_R input1 (.A(enable_i),
    .Y(net2));
 BUFx2_ASAP7_75t_R output2 (.A(net21),
    .Y(counter_value_o[0]));
 BUFx2_ASAP7_75t_R output3 (.A(net25),
    .Y(counter_value_o[1]));
 BUFx3_ASAP7_75t_R output4 (.A(net5),
    .Y(counter_value_o[2]));
 BUFx3_ASAP7_75t_R output5 (.A(net6),
    .Y(counter_value_o[3]));
 TIEHIx1_ASAP7_75t_R \counter_0.n20_q[0]$_DFFE_PN0P__6  (.H(net7));
 TIEHIx1_ASAP7_75t_R \counter_0.n20_q[1]$_DFFE_PN0P__7  (.H(net8));
 TIEHIx1_ASAP7_75t_R \counter_0.n20_q[2]$_DFFE_PN0P__8  (.H(net9));
 TIEHIx1_ASAP7_75t_R \counter_0.n20_q[3]$_DFFE_PN0P__9  (.H(net10));
 BUFx2_ASAP7_75t_R clkbuf_1_0__f_clock_i (.A(clknet_0_clock_i),
    .Y(clknet_1_0__leaf_clock_i));
 BUFx2_ASAP7_75t_R clkbuf_1_1__f_clock_i (.A(clknet_0_clock_i),
    .Y(clknet_1_1__leaf_clock_i));
 BUFx3_ASAP7_75t_R rebuffer1 (.A(_04_),
    .Y(net11));
 BUFx3_ASAP7_75t_R rebuffer2 (.A(_04_),
    .Y(net12));
 BUFx2_ASAP7_75t_R rebuffer3 (.A(net17),
    .Y(net13));
 BUFx2_ASAP7_75t_R rebuffer4 (.A(net26),
    .Y(net14));
 BUFx2_ASAP7_75t_R rebuffer5 (.A(_02_),
    .Y(net15));
 BUFx2_ASAP7_75t_R rebuffer6 (.A(net19),
    .Y(net16));
 BUFx2_ASAP7_75t_R rebuffer7 (.A(net18),
    .Y(net17));
 BUFx2_ASAP7_75t_R rebuffer8 (.A(_03_),
    .Y(net18));
 BUFx2_ASAP7_75t_R rebuffer9 (.A(net20),
    .Y(net19));
 BUFx2_ASAP7_75t_R rebuffer10 (.A(_02_),
    .Y(net20));
 BUFx2_ASAP7_75t_R rebuffer11 (.A(net3),
    .Y(net21));
 BUFx2_ASAP7_75t_R rebuffer12 (.A(_01_),
    .Y(net22));
 BUFx3_ASAP7_75t_R rebuffer13 (.A(_01_),
    .Y(net23));
 BUFx2_ASAP7_75t_R hold14 (.A(reset_n_i),
    .Y(net24));
 BUFx2_ASAP7_75t_R rebuffer14 (.A(net4),
    .Y(net25));
 BUFx2_ASAP7_75t_R rebuffer15 (.A(_03_),
    .Y(net26));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx4_ASAP7_75t_R FILLER_1_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_144 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx4_ASAP7_75t_R FILLER_2_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_144 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx4_ASAP7_75t_R FILLER_3_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_144 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_4_112 ();
 DECAPx4_ASAP7_75t_R FILLER_4_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_144 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_5_112 ();
 DECAPx4_ASAP7_75t_R FILLER_5_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_144 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_6_112 ();
 DECAPx4_ASAP7_75t_R FILLER_6_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_144 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_7_112 ();
 DECAPx4_ASAP7_75t_R FILLER_7_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_144 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_8_112 ();
 DECAPx4_ASAP7_75t_R FILLER_8_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_144 ();
 DECAPx2_ASAP7_75t_R FILLER_9_2 ();
 FILLER_ASAP7_75t_R FILLER_9_8 ();
 DECAPx10_ASAP7_75t_R FILLER_9_15 ();
 DECAPx10_ASAP7_75t_R FILLER_9_37 ();
 DECAPx10_ASAP7_75t_R FILLER_9_59 ();
 DECAPx10_ASAP7_75t_R FILLER_9_81 ();
 DECAPx10_ASAP7_75t_R FILLER_9_103 ();
 DECAPx6_ASAP7_75t_R FILLER_9_125 ();
 DECAPx2_ASAP7_75t_R FILLER_9_139 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_112 ();
 DECAPx4_ASAP7_75t_R FILLER_10_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_144 ();
 DECAPx2_ASAP7_75t_R FILLER_11_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_14 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_27 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_33 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_38 ();
 DECAPx10_ASAP7_75t_R FILLER_11_49 ();
 DECAPx10_ASAP7_75t_R FILLER_11_71 ();
 DECAPx10_ASAP7_75t_R FILLER_11_93 ();
 DECAPx10_ASAP7_75t_R FILLER_11_115 ();
 DECAPx2_ASAP7_75t_R FILLER_11_137 ();
 FILLER_ASAP7_75t_R FILLER_11_143 ();
 FILLER_ASAP7_75t_R FILLER_12_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_30 ();
 FILLER_ASAP7_75t_R FILLER_12_37 ();
 DECAPx10_ASAP7_75t_R FILLER_12_60 ();
 DECAPx10_ASAP7_75t_R FILLER_12_82 ();
 DECAPx10_ASAP7_75t_R FILLER_12_104 ();
 DECAPx6_ASAP7_75t_R FILLER_12_126 ();
 DECAPx1_ASAP7_75t_R FILLER_12_140 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_2 ();
 FILLER_ASAP7_75t_R FILLER_13_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_36 ();
 DECAPx10_ASAP7_75t_R FILLER_13_67 ();
 DECAPx10_ASAP7_75t_R FILLER_13_89 ();
 DECAPx10_ASAP7_75t_R FILLER_13_111 ();
 DECAPx4_ASAP7_75t_R FILLER_13_133 ();
 FILLER_ASAP7_75t_R FILLER_13_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_48 ();
 DECAPx10_ASAP7_75t_R FILLER_14_71 ();
 DECAPx10_ASAP7_75t_R FILLER_14_93 ();
 DECAPx10_ASAP7_75t_R FILLER_14_115 ();
 DECAPx2_ASAP7_75t_R FILLER_14_137 ();
 FILLER_ASAP7_75t_R FILLER_14_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_8 ();
 DECAPx10_ASAP7_75t_R FILLER_15_63 ();
 DECAPx4_ASAP7_75t_R FILLER_15_85 ();
 FILLER_ASAP7_75t_R FILLER_15_95 ();
 DECAPx10_ASAP7_75t_R FILLER_15_102 ();
 DECAPx6_ASAP7_75t_R FILLER_15_124 ();
 DECAPx2_ASAP7_75t_R FILLER_15_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_144 ();
 DECAPx1_ASAP7_75t_R FILLER_16_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_6 ();
 FILLER_ASAP7_75t_R FILLER_16_12 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_14 ();
 FILLER_ASAP7_75t_R FILLER_16_20 ();
 DECAPx10_ASAP7_75t_R FILLER_16_59 ();
 DECAPx10_ASAP7_75t_R FILLER_16_81 ();
 DECAPx10_ASAP7_75t_R FILLER_16_103 ();
 DECAPx6_ASAP7_75t_R FILLER_16_125 ();
 DECAPx2_ASAP7_75t_R FILLER_16_139 ();
 DECAPx6_ASAP7_75t_R FILLER_17_2 ();
 DECAPx1_ASAP7_75t_R FILLER_17_16 ();
 DECAPx2_ASAP7_75t_R FILLER_17_23 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_29 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_34 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_40 ();
 DECAPx10_ASAP7_75t_R FILLER_17_46 ();
 DECAPx10_ASAP7_75t_R FILLER_17_68 ();
 DECAPx10_ASAP7_75t_R FILLER_17_90 ();
 DECAPx10_ASAP7_75t_R FILLER_17_112 ();
 DECAPx4_ASAP7_75t_R FILLER_17_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_144 ();
 DECAPx10_ASAP7_75t_R FILLER_18_2 ();
 DECAPx10_ASAP7_75t_R FILLER_18_24 ();
 DECAPx10_ASAP7_75t_R FILLER_18_46 ();
 DECAPx10_ASAP7_75t_R FILLER_18_68 ();
 DECAPx10_ASAP7_75t_R FILLER_18_90 ();
 DECAPx10_ASAP7_75t_R FILLER_18_112 ();
 DECAPx4_ASAP7_75t_R FILLER_18_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_144 ();
 DECAPx1_ASAP7_75t_R FILLER_19_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_6 ();
 DECAPx10_ASAP7_75t_R FILLER_19_12 ();
 DECAPx10_ASAP7_75t_R FILLER_19_34 ();
 DECAPx10_ASAP7_75t_R FILLER_19_56 ();
 DECAPx10_ASAP7_75t_R FILLER_19_78 ();
 DECAPx10_ASAP7_75t_R FILLER_19_100 ();
 DECAPx10_ASAP7_75t_R FILLER_19_122 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_144 ();
 DECAPx10_ASAP7_75t_R FILLER_20_2 ();
 DECAPx10_ASAP7_75t_R FILLER_20_24 ();
 DECAPx10_ASAP7_75t_R FILLER_20_46 ();
 DECAPx10_ASAP7_75t_R FILLER_20_68 ();
 DECAPx10_ASAP7_75t_R FILLER_20_90 ();
 DECAPx10_ASAP7_75t_R FILLER_20_112 ();
 DECAPx4_ASAP7_75t_R FILLER_20_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_20_144 ();
 DECAPx10_ASAP7_75t_R FILLER_21_2 ();
 DECAPx10_ASAP7_75t_R FILLER_21_24 ();
 DECAPx10_ASAP7_75t_R FILLER_21_46 ();
 DECAPx10_ASAP7_75t_R FILLER_21_68 ();
 DECAPx10_ASAP7_75t_R FILLER_21_90 ();
 DECAPx10_ASAP7_75t_R FILLER_21_112 ();
 DECAPx4_ASAP7_75t_R FILLER_21_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_144 ();
 DECAPx10_ASAP7_75t_R FILLER_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_22_68 ();
 DECAPx10_ASAP7_75t_R FILLER_22_90 ();
 DECAPx10_ASAP7_75t_R FILLER_22_112 ();
 DECAPx4_ASAP7_75t_R FILLER_22_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_144 ();
 DECAPx10_ASAP7_75t_R FILLER_23_2 ();
 DECAPx10_ASAP7_75t_R FILLER_23_24 ();
 DECAPx10_ASAP7_75t_R FILLER_23_46 ();
 DECAPx10_ASAP7_75t_R FILLER_23_68 ();
 DECAPx10_ASAP7_75t_R FILLER_23_90 ();
 DECAPx10_ASAP7_75t_R FILLER_23_112 ();
 DECAPx4_ASAP7_75t_R FILLER_23_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_23_144 ();
 DECAPx10_ASAP7_75t_R FILLER_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_24_68 ();
 DECAPx10_ASAP7_75t_R FILLER_24_90 ();
 DECAPx10_ASAP7_75t_R FILLER_24_112 ();
 DECAPx4_ASAP7_75t_R FILLER_24_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_144 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_25_68 ();
 DECAPx10_ASAP7_75t_R FILLER_25_90 ();
 DECAPx10_ASAP7_75t_R FILLER_25_112 ();
 DECAPx4_ASAP7_75t_R FILLER_25_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_144 ();
 DECAPx10_ASAP7_75t_R FILLER_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_26_68 ();
 DECAPx10_ASAP7_75t_R FILLER_26_90 ();
 DECAPx10_ASAP7_75t_R FILLER_26_112 ();
 DECAPx4_ASAP7_75t_R FILLER_26_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_144 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_27_46 ();
 DECAPx10_ASAP7_75t_R FILLER_27_68 ();
 DECAPx10_ASAP7_75t_R FILLER_27_90 ();
 DECAPx10_ASAP7_75t_R FILLER_27_112 ();
 DECAPx4_ASAP7_75t_R FILLER_27_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_144 ();
 DECAPx10_ASAP7_75t_R FILLER_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_28_46 ();
 DECAPx10_ASAP7_75t_R FILLER_28_68 ();
 DECAPx10_ASAP7_75t_R FILLER_28_90 ();
 DECAPx10_ASAP7_75t_R FILLER_28_112 ();
 DECAPx4_ASAP7_75t_R FILLER_28_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_144 ();
endmodule
