module counter_board (clock_i,
    enable_i,
    reset_n_i,
    counter_value_o);
 input clock_i;
 input enable_i;
 input reset_n_i;
 output [3:0] counter_value_o;

 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire n1_o;
 wire \counter_0/_00_ ;
 wire \counter_0/_01_ ;
 wire \counter_0/_02_ ;
 wire \counter_0/_03_ ;
 wire \counter_0/_04_ ;
 wire \counter_0/_05_ ;
 wire \counter_0/_06_ ;
 wire \counter_0/_07_ ;
 wire \counter_0/_08_ ;
 wire \counter_0/_09_ ;
 wire \counter_0/_10_ ;
 wire \counter_0/_11_ ;
 wire \counter_0/_12_ ;
 wire \counter_0/_13_ ;
 wire \counter_0/_14_ ;
 wire \counter_0/_15_ ;
 wire \counter_0/_16_ ;
 wire \counter_0/_17_ ;
 wire \counter_0/_18_ ;
 wire clknet_0_clock_i;
 wire net1;
 wire net2;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire clknet_1_0__leaf_clock_i;
 wire clknet_1_1__leaf_clock_i;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net19;

 INVx3_ASAP7_75t_R _0_ (.A(net2),
    .Y(n1_o));
 INVx2_ASAP7_75t_R \counter_0/_20_  (.A(\counter_0/_01_ ),
    .Y(net5));
 INVx1_ASAP7_75t_R \counter_0/_21_  (.A(\counter_0/_00_ ),
    .Y(net6));
 INVx2_ASAP7_75t_R \counter_0/_22_  (.A(\counter_0/_02_ ),
    .Y(net4));
 INVx2_ASAP7_75t_R \counter_0/_23_  (.A(\counter_0/_03_ ),
    .Y(net3));
 INVx2_ASAP7_75t_R \counter_0/_24_  (.A(n1_o),
    .Y(\counter_0/_06_ ));
 INVx2_ASAP7_75t_R \counter_0/_25_  (.A(net1),
    .Y(\counter_0/_11_ ));
 OR3x1_ASAP7_75t_R \counter_0/_26_  (.A(\counter_0/_04_ ),
    .B(\counter_0/_01_ ),
    .C(\counter_0/_00_ ),
    .Y(\counter_0/_12_ ));
 AND3x1_ASAP7_75t_R \counter_0/_27_  (.A(\counter_0/_12_ ),
    .B(net1),
    .C(net14),
    .Y(\counter_0/_13_ ));
 AO21x1_ASAP7_75t_R \counter_0/_28_  (.A1(net3),
    .A2(\counter_0/_11_ ),
    .B(\counter_0/_13_ ),
    .Y(\counter_0/_07_ ));
 NAND2x1_ASAP7_75t_R \counter_0/_29_  (.A(net1),
    .B(\counter_0/_05_ ),
    .Y(\counter_0/_14_ ));
 OA21x2_ASAP7_75t_R \counter_0/_30_  (.A1(net18),
    .A2(net1),
    .B(\counter_0/_14_ ),
    .Y(\counter_0/_08_ ));
 NOR2x2_ASAP7_75t_R \counter_0/_31_  (.A(net11),
    .B(\counter_0/_11_ ),
    .Y(\counter_0/_15_ ));
 XNOR2x1_ASAP7_75t_R \counter_0/_32_  (.B(\counter_0/_15_ ),
    .Y(\counter_0/_09_ ),
    .A(net25));
 OR4x1_ASAP7_75t_R \counter_0/_33_  (.A(\counter_0/_01_ ),
    .B(net15),
    .C(\counter_0/_03_ ),
    .D(\counter_0/_11_ ),
    .Y(\counter_0/_16_ ));
 OAI21x1_ASAP7_75t_R \counter_0/_34_  (.A1(net19),
    .A2(net13),
    .B(net12),
    .Y(\counter_0/_17_ ));
 AND4x1_ASAP7_75t_R \counter_0/_35_  (.A(\counter_0/_17_ ),
    .B(net5),
    .C(net1),
    .D(net6),
    .Y(\counter_0/_18_ ));
 AOI21x1_ASAP7_75t_R \counter_0/_36_  (.A1(\counter_0/_00_ ),
    .A2(\counter_0/_16_ ),
    .B(\counter_0/_18_ ),
    .Y(\counter_0/_10_ ));
 HAxp5_ASAP7_75t_R \counter_0/_37_  (.A(net3),
    .B(net4),
    .CON(\counter_0/_04_ ),
    .SN(\counter_0/_05_ ));
 BUFx2_ASAP7_75t_R clkbuf_0_clock_i (.A(clock_i),
    .Y(clknet_0_clock_i));
 DFFASRHQNx1_ASAP7_75t_R \counter_0/n20_q[0]$_DFFE_PP0P_  (.CLK(clknet_1_0__leaf_clock_i),
    .D(\counter_0/_07_ ),
    .QN(\counter_0/_03_ ),
    .RESETN(net7),
    .SETN(\counter_0/_06_ ));
 DFFASRHQNx1_ASAP7_75t_R \counter_0/n20_q[1]$_DFFE_PP0P_  (.CLK(clknet_1_0__leaf_clock_i),
    .D(\counter_0/_08_ ),
    .QN(\counter_0/_02_ ),
    .RESETN(net8),
    .SETN(\counter_0/_06_ ));
 DFFASRHQNx1_ASAP7_75t_R \counter_0/n20_q[2]$_DFFE_PP0P_  (.CLK(clknet_1_1__leaf_clock_i),
    .D(\counter_0/_09_ ),
    .QN(\counter_0/_01_ ),
    .RESETN(net9),
    .SETN(\counter_0/_06_ ));
 DFFASRHQNx1_ASAP7_75t_R \counter_0/n20_q[3]$_DFFE_PP0P_  (.CLK(clknet_1_1__leaf_clock_i),
    .D(\counter_0/_10_ ),
    .QN(\counter_0/_00_ ),
    .RESETN(net10),
    .SETN(\counter_0/_06_ ));
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Right_0 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Right_1 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Right_2 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Right_3 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Right_4 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Right_5 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Right_6 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Right_7 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Right_8 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Right_9 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Right_10 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Right_11 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Right_12 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Right_13 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Right_14 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Right_15 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Right_16 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Right_17 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Right_18 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Right_19 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Right_20 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Right_21 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Right_22 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Right_23 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Right_24 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Right_25 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Right_26 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Right_27 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Right_28 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_0_Left_29 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_1_Left_30 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_2_Left_31 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_3_Left_32 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_4_Left_33 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_5_Left_34 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_6_Left_35 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_7_Left_36 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_8_Left_37 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_9_Left_38 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_10_Left_39 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_11_Left_40 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_12_Left_41 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_13_Left_42 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_14_Left_43 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_15_Left_44 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_16_Left_45 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_17_Left_46 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_18_Left_47 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_19_Left_48 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_20_Left_49 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_21_Left_50 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_22_Left_51 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_23_Left_52 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_24_Left_53 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_25_Left_54 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_26_Left_55 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_27_Left_56 ();
 TAPCELL_ASAP7_75t_R PHY_EDGE_ROW_28_Left_57 ();
 BUFx2_ASAP7_75t_R input1 (.A(enable_i),
    .Y(net1));
 BUFx2_ASAP7_75t_R input2 (.A(reset_n_i),
    .Y(net2));
 BUFx2_ASAP7_75t_R output3 (.A(net24),
    .Y(counter_value_o[0]));
 BUFx3_ASAP7_75t_R output4 (.A(net18),
    .Y(counter_value_o[1]));
 BUFx2_ASAP7_75t_R output5 (.A(net5),
    .Y(counter_value_o[2]));
 BUFx3_ASAP7_75t_R output6 (.A(net6),
    .Y(counter_value_o[3]));
 TIEHIx1_ASAP7_75t_R \counter_0/n20_q[0]$_DFFE_PP0P__7  (.H(net7));
 TIEHIx1_ASAP7_75t_R \counter_0/n20_q[1]$_DFFE_PP0P__8  (.H(net8));
 TIEHIx1_ASAP7_75t_R \counter_0/n20_q[2]$_DFFE_PP0P__9  (.H(net9));
 TIEHIx1_ASAP7_75t_R \counter_0/n20_q[3]$_DFFE_PP0P__10  (.H(net10));
 BUFx2_ASAP7_75t_R clkbuf_1_0__f_clock_i (.A(clknet_0_clock_i),
    .Y(clknet_1_0__leaf_clock_i));
 BUFx2_ASAP7_75t_R clkbuf_1_1__f_clock_i (.A(clknet_0_clock_i),
    .Y(clknet_1_1__leaf_clock_i));
 BUFx3_ASAP7_75t_R rebuffer1 (.A(\counter_0/_04_ ),
    .Y(net11));
 BUFx3_ASAP7_75t_R rebuffer2 (.A(\counter_0/_04_ ),
    .Y(net12));
 BUFx2_ASAP7_75t_R rebuffer3 (.A(\counter_0/_03_ ),
    .Y(net13));
 BUFx2_ASAP7_75t_R rebuffer4 (.A(net22),
    .Y(net14));
 BUFx3_ASAP7_75t_R rebuffer5 (.A(net16),
    .Y(net15));
 BUFx3_ASAP7_75t_R rebuffer6 (.A(net17),
    .Y(net16));
 BUFx3_ASAP7_75t_R rebuffer7 (.A(\counter_0/_02_ ),
    .Y(net17));
 BUFx3_ASAP7_75t_R rebuffer8 (.A(net4),
    .Y(net18));
 BUFx2_ASAP7_75t_R rebuffer12 (.A(net23),
    .Y(net22));
 BUFx2_ASAP7_75t_R rebuffer13 (.A(\counter_0/_03_ ),
    .Y(net23));
 BUFx2_ASAP7_75t_R rebuffer14 (.A(net3),
    .Y(net24));
 BUFx2_ASAP7_75t_R rebuffer15 (.A(\counter_0/_01_ ),
    .Y(net25));
 BUFx2_ASAP7_75t_R rebuffer9 (.A(\counter_0/_02_ ),
    .Y(net19));
 DECAPx10_ASAP7_75t_R FILLER_0_2 ();
 DECAPx10_ASAP7_75t_R FILLER_0_24 ();
 DECAPx10_ASAP7_75t_R FILLER_0_46 ();
 DECAPx10_ASAP7_75t_R FILLER_0_68 ();
 DECAPx10_ASAP7_75t_R FILLER_0_90 ();
 DECAPx10_ASAP7_75t_R FILLER_0_112 ();
 DECAPx4_ASAP7_75t_R FILLER_0_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_0_144 ();
 DECAPx10_ASAP7_75t_R FILLER_1_2 ();
 DECAPx10_ASAP7_75t_R FILLER_1_24 ();
 DECAPx10_ASAP7_75t_R FILLER_1_46 ();
 DECAPx10_ASAP7_75t_R FILLER_1_68 ();
 DECAPx10_ASAP7_75t_R FILLER_1_90 ();
 DECAPx10_ASAP7_75t_R FILLER_1_112 ();
 DECAPx4_ASAP7_75t_R FILLER_1_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_1_144 ();
 DECAPx10_ASAP7_75t_R FILLER_2_2 ();
 DECAPx10_ASAP7_75t_R FILLER_2_24 ();
 DECAPx10_ASAP7_75t_R FILLER_2_46 ();
 DECAPx10_ASAP7_75t_R FILLER_2_68 ();
 DECAPx10_ASAP7_75t_R FILLER_2_90 ();
 DECAPx10_ASAP7_75t_R FILLER_2_112 ();
 DECAPx4_ASAP7_75t_R FILLER_2_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_2_144 ();
 DECAPx10_ASAP7_75t_R FILLER_3_2 ();
 DECAPx10_ASAP7_75t_R FILLER_3_24 ();
 DECAPx10_ASAP7_75t_R FILLER_3_46 ();
 DECAPx10_ASAP7_75t_R FILLER_3_68 ();
 DECAPx10_ASAP7_75t_R FILLER_3_90 ();
 DECAPx10_ASAP7_75t_R FILLER_3_112 ();
 DECAPx4_ASAP7_75t_R FILLER_3_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_3_144 ();
 DECAPx10_ASAP7_75t_R FILLER_4_2 ();
 DECAPx10_ASAP7_75t_R FILLER_4_24 ();
 DECAPx10_ASAP7_75t_R FILLER_4_46 ();
 DECAPx10_ASAP7_75t_R FILLER_4_68 ();
 DECAPx10_ASAP7_75t_R FILLER_4_90 ();
 DECAPx10_ASAP7_75t_R FILLER_4_112 ();
 DECAPx4_ASAP7_75t_R FILLER_4_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_4_144 ();
 DECAPx10_ASAP7_75t_R FILLER_5_2 ();
 DECAPx10_ASAP7_75t_R FILLER_5_24 ();
 DECAPx10_ASAP7_75t_R FILLER_5_46 ();
 DECAPx10_ASAP7_75t_R FILLER_5_68 ();
 DECAPx10_ASAP7_75t_R FILLER_5_90 ();
 DECAPx10_ASAP7_75t_R FILLER_5_112 ();
 DECAPx4_ASAP7_75t_R FILLER_5_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_5_144 ();
 DECAPx10_ASAP7_75t_R FILLER_6_2 ();
 DECAPx10_ASAP7_75t_R FILLER_6_24 ();
 DECAPx10_ASAP7_75t_R FILLER_6_46 ();
 DECAPx10_ASAP7_75t_R FILLER_6_68 ();
 DECAPx10_ASAP7_75t_R FILLER_6_90 ();
 DECAPx10_ASAP7_75t_R FILLER_6_112 ();
 DECAPx4_ASAP7_75t_R FILLER_6_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_6_144 ();
 DECAPx10_ASAP7_75t_R FILLER_7_2 ();
 DECAPx10_ASAP7_75t_R FILLER_7_24 ();
 DECAPx10_ASAP7_75t_R FILLER_7_46 ();
 DECAPx10_ASAP7_75t_R FILLER_7_68 ();
 DECAPx10_ASAP7_75t_R FILLER_7_90 ();
 DECAPx10_ASAP7_75t_R FILLER_7_112 ();
 DECAPx4_ASAP7_75t_R FILLER_7_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_7_144 ();
 DECAPx10_ASAP7_75t_R FILLER_8_2 ();
 DECAPx10_ASAP7_75t_R FILLER_8_24 ();
 DECAPx10_ASAP7_75t_R FILLER_8_46 ();
 DECAPx10_ASAP7_75t_R FILLER_8_68 ();
 DECAPx10_ASAP7_75t_R FILLER_8_90 ();
 DECAPx10_ASAP7_75t_R FILLER_8_112 ();
 DECAPx4_ASAP7_75t_R FILLER_8_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_8_144 ();
 DECAPx10_ASAP7_75t_R FILLER_9_2 ();
 DECAPx10_ASAP7_75t_R FILLER_9_24 ();
 DECAPx10_ASAP7_75t_R FILLER_9_46 ();
 DECAPx10_ASAP7_75t_R FILLER_9_68 ();
 DECAPx10_ASAP7_75t_R FILLER_9_90 ();
 DECAPx10_ASAP7_75t_R FILLER_9_112 ();
 DECAPx4_ASAP7_75t_R FILLER_9_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_9_144 ();
 DECAPx10_ASAP7_75t_R FILLER_10_2 ();
 DECAPx10_ASAP7_75t_R FILLER_10_24 ();
 DECAPx10_ASAP7_75t_R FILLER_10_46 ();
 DECAPx10_ASAP7_75t_R FILLER_10_68 ();
 DECAPx10_ASAP7_75t_R FILLER_10_90 ();
 DECAPx10_ASAP7_75t_R FILLER_10_112 ();
 DECAPx4_ASAP7_75t_R FILLER_10_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_10_144 ();
 DECAPx10_ASAP7_75t_R FILLER_11_2 ();
 DECAPx10_ASAP7_75t_R FILLER_11_24 ();
 DECAPx10_ASAP7_75t_R FILLER_11_46 ();
 DECAPx10_ASAP7_75t_R FILLER_11_68 ();
 DECAPx10_ASAP7_75t_R FILLER_11_90 ();
 DECAPx10_ASAP7_75t_R FILLER_11_112 ();
 DECAPx4_ASAP7_75t_R FILLER_11_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_11_144 ();
 DECAPx10_ASAP7_75t_R FILLER_12_2 ();
 DECAPx10_ASAP7_75t_R FILLER_12_24 ();
 DECAPx10_ASAP7_75t_R FILLER_12_46 ();
 DECAPx10_ASAP7_75t_R FILLER_12_68 ();
 DECAPx10_ASAP7_75t_R FILLER_12_90 ();
 DECAPx10_ASAP7_75t_R FILLER_12_112 ();
 DECAPx4_ASAP7_75t_R FILLER_12_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_12_144 ();
 DECAPx10_ASAP7_75t_R FILLER_13_2 ();
 DECAPx10_ASAP7_75t_R FILLER_13_24 ();
 DECAPx10_ASAP7_75t_R FILLER_13_46 ();
 DECAPx10_ASAP7_75t_R FILLER_13_68 ();
 DECAPx10_ASAP7_75t_R FILLER_13_90 ();
 DECAPx10_ASAP7_75t_R FILLER_13_112 ();
 DECAPx4_ASAP7_75t_R FILLER_13_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_13_144 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_2 ();
 FILLER_ASAP7_75t_R FILLER_14_9 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_11 ();
 DECAPx10_ASAP7_75t_R FILLER_14_28 ();
 DECAPx10_ASAP7_75t_R FILLER_14_50 ();
 DECAPx10_ASAP7_75t_R FILLER_14_72 ();
 DECAPx10_ASAP7_75t_R FILLER_14_94 ();
 DECAPx10_ASAP7_75t_R FILLER_14_116 ();
 DECAPx2_ASAP7_75t_R FILLER_14_138 ();
 FILLERxp5_ASAP7_75t_R FILLER_14_144 ();
 DECAPx6_ASAP7_75t_R FILLER_15_2 ();
 DECAPx2_ASAP7_75t_R FILLER_15_16 ();
 FILLERxp5_ASAP7_75t_R FILLER_15_22 ();
 DECAPx2_ASAP7_75t_R FILLER_15_28 ();
 FILLER_ASAP7_75t_R FILLER_15_34 ();
 DECAPx10_ASAP7_75t_R FILLER_15_41 ();
 DECAPx10_ASAP7_75t_R FILLER_15_63 ();
 DECAPx10_ASAP7_75t_R FILLER_15_85 ();
 DECAPx10_ASAP7_75t_R FILLER_15_107 ();
 DECAPx6_ASAP7_75t_R FILLER_15_129 ();
 FILLER_ASAP7_75t_R FILLER_15_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_16_2 ();
 DECAPx10_ASAP7_75t_R FILLER_16_60 ();
 DECAPx10_ASAP7_75t_R FILLER_16_82 ();
 DECAPx10_ASAP7_75t_R FILLER_16_104 ();
 DECAPx2_ASAP7_75t_R FILLER_16_126 ();
 DECAPx2_ASAP7_75t_R FILLER_16_137 ();
 FILLER_ASAP7_75t_R FILLER_16_143 ();
 DECAPx2_ASAP7_75t_R FILLER_17_2 ();
 FILLER_ASAP7_75t_R FILLER_17_8 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_10 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_54 ();
 DECAPx10_ASAP7_75t_R FILLER_17_66 ();
 DECAPx10_ASAP7_75t_R FILLER_17_88 ();
 DECAPx10_ASAP7_75t_R FILLER_17_110 ();
 DECAPx4_ASAP7_75t_R FILLER_17_132 ();
 FILLER_ASAP7_75t_R FILLER_17_142 ();
 FILLERxp5_ASAP7_75t_R FILLER_17_144 ();
 FILLER_ASAP7_75t_R FILLER_18_2 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_4 ();
 FILLER_ASAP7_75t_R FILLER_18_39 ();
 FILLERxp5_ASAP7_75t_R FILLER_18_41 ();
 DECAPx10_ASAP7_75t_R FILLER_18_67 ();
 DECAPx10_ASAP7_75t_R FILLER_18_89 ();
 DECAPx10_ASAP7_75t_R FILLER_18_111 ();
 DECAPx4_ASAP7_75t_R FILLER_18_133 ();
 FILLER_ASAP7_75t_R FILLER_18_143 ();
 FILLERxp5_ASAP7_75t_R FILLER_19_2 ();
 FILLER_ASAP7_75t_R FILLER_19_29 ();
 DECAPx10_ASAP7_75t_R FILLER_19_71 ();
 DECAPx10_ASAP7_75t_R FILLER_19_93 ();
 DECAPx10_ASAP7_75t_R FILLER_19_115 ();
 DECAPx2_ASAP7_75t_R FILLER_19_137 ();
 FILLER_ASAP7_75t_R FILLER_19_143 ();
 DECAPx2_ASAP7_75t_R FILLER_20_2 ();
 FILLER_ASAP7_75t_R FILLER_20_20 ();
 FILLER_ASAP7_75t_R FILLER_20_32 ();
 DECAPx10_ASAP7_75t_R FILLER_20_65 ();
 DECAPx10_ASAP7_75t_R FILLER_20_87 ();
 DECAPx10_ASAP7_75t_R FILLER_20_109 ();
 DECAPx6_ASAP7_75t_R FILLER_20_131 ();
 DECAPx6_ASAP7_75t_R FILLER_21_2 ();
 DECAPx2_ASAP7_75t_R FILLER_21_16 ();
 DECAPx1_ASAP7_75t_R FILLER_21_25 ();
 DECAPx2_ASAP7_75t_R FILLER_21_34 ();
 FILLER_ASAP7_75t_R FILLER_21_40 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_42 ();
 FILLER_ASAP7_75t_R FILLER_21_48 ();
 FILLERxp5_ASAP7_75t_R FILLER_21_50 ();
 DECAPx10_ASAP7_75t_R FILLER_21_61 ();
 DECAPx10_ASAP7_75t_R FILLER_21_83 ();
 DECAPx10_ASAP7_75t_R FILLER_21_105 ();
 DECAPx6_ASAP7_75t_R FILLER_21_127 ();
 DECAPx1_ASAP7_75t_R FILLER_21_141 ();
 DECAPx10_ASAP7_75t_R FILLER_22_2 ();
 DECAPx10_ASAP7_75t_R FILLER_22_24 ();
 DECAPx10_ASAP7_75t_R FILLER_22_46 ();
 DECAPx10_ASAP7_75t_R FILLER_22_68 ();
 DECAPx10_ASAP7_75t_R FILLER_22_90 ();
 DECAPx10_ASAP7_75t_R FILLER_22_112 ();
 DECAPx4_ASAP7_75t_R FILLER_22_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_22_144 ();
 DECAPx2_ASAP7_75t_R FILLER_23_2 ();
 FILLER_ASAP7_75t_R FILLER_23_8 ();
 DECAPx10_ASAP7_75t_R FILLER_23_15 ();
 DECAPx10_ASAP7_75t_R FILLER_23_37 ();
 DECAPx10_ASAP7_75t_R FILLER_23_59 ();
 DECAPx10_ASAP7_75t_R FILLER_23_81 ();
 DECAPx10_ASAP7_75t_R FILLER_23_103 ();
 DECAPx6_ASAP7_75t_R FILLER_23_125 ();
 DECAPx2_ASAP7_75t_R FILLER_23_139 ();
 DECAPx10_ASAP7_75t_R FILLER_24_2 ();
 DECAPx10_ASAP7_75t_R FILLER_24_24 ();
 DECAPx10_ASAP7_75t_R FILLER_24_46 ();
 DECAPx10_ASAP7_75t_R FILLER_24_68 ();
 DECAPx10_ASAP7_75t_R FILLER_24_90 ();
 DECAPx10_ASAP7_75t_R FILLER_24_112 ();
 DECAPx4_ASAP7_75t_R FILLER_24_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_24_144 ();
 DECAPx10_ASAP7_75t_R FILLER_25_2 ();
 DECAPx10_ASAP7_75t_R FILLER_25_24 ();
 DECAPx10_ASAP7_75t_R FILLER_25_46 ();
 DECAPx10_ASAP7_75t_R FILLER_25_68 ();
 DECAPx10_ASAP7_75t_R FILLER_25_90 ();
 DECAPx10_ASAP7_75t_R FILLER_25_112 ();
 DECAPx4_ASAP7_75t_R FILLER_25_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_25_144 ();
 DECAPx10_ASAP7_75t_R FILLER_26_2 ();
 DECAPx10_ASAP7_75t_R FILLER_26_24 ();
 DECAPx10_ASAP7_75t_R FILLER_26_46 ();
 DECAPx10_ASAP7_75t_R FILLER_26_68 ();
 DECAPx10_ASAP7_75t_R FILLER_26_90 ();
 DECAPx10_ASAP7_75t_R FILLER_26_112 ();
 DECAPx4_ASAP7_75t_R FILLER_26_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_26_144 ();
 DECAPx10_ASAP7_75t_R FILLER_27_2 ();
 DECAPx10_ASAP7_75t_R FILLER_27_24 ();
 DECAPx10_ASAP7_75t_R FILLER_27_46 ();
 DECAPx10_ASAP7_75t_R FILLER_27_68 ();
 DECAPx10_ASAP7_75t_R FILLER_27_90 ();
 DECAPx10_ASAP7_75t_R FILLER_27_112 ();
 DECAPx4_ASAP7_75t_R FILLER_27_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_27_144 ();
 DECAPx10_ASAP7_75t_R FILLER_28_2 ();
 DECAPx10_ASAP7_75t_R FILLER_28_24 ();
 DECAPx10_ASAP7_75t_R FILLER_28_46 ();
 DECAPx10_ASAP7_75t_R FILLER_28_68 ();
 DECAPx10_ASAP7_75t_R FILLER_28_90 ();
 DECAPx10_ASAP7_75t_R FILLER_28_112 ();
 DECAPx4_ASAP7_75t_R FILLER_28_134 ();
 FILLERxp5_ASAP7_75t_R FILLER_28_144 ();
endmodule
